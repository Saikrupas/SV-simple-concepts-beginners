/*

Assignment 4:-  Generate 25 stimuli for the Code mentioned in Instruction tab

Refer methodology discussed in the previous lecture and 
try to generate 25 stimuli for testing the system mentioned in the Instruction Tab.

Generate 25 stimuli for the code mentioned below. Use methodology 
discussed in the previous lecture. Use of the Generator and Driver is prohibited.

Try to add for loop in the Testbench top to apply 25 stimuli to DUT. 
Stimulus generation will happen in the Testbench top. 
Your task should be to capture the response of DUT in Monitor as well as Scoreboard.

Refer snippets --> Assignment-4(Section-6) snippet, Assignment-4(Section-6) snippet-2
*/